/*
   CS/ECE 552 Spring '20
  
   Filename        : decode.v
   Description     : This is the module for the overall decode stage of the processor.
*/
module decode (/* TODO: Add appropriate inputs/outputs for your decode stage here*/);

   // TODO: Your code here
   
endmodule
