/*
   CS/ECE 552 Spring '20
  
   Filename        : fetch.v
   Description     : This is the module for the overall fetch stage of the processor.
*/
module fetch (clk, rst, /*err,*/ stall, 
               branch_jump_pc, PCSrc, Jump_IDEX,
               Halt_fetch, pcAdd2, 
               inst_mem_err,
               inst_mem_stall,
               inst_mem_done,
               instruction
               );
   /* TODO: Add appropriate inputs/outputs for your fetch stage here*/
   
   input clk,rst;
   input stall;
   input [15:0] branch_jump_pc;  //used to be next_pc2
   input PCSrc;                  //branch_jump_taken signal
   input Jump_IDEX;
   input Halt_fetch;
   output [15:0] pcAdd2; //PC+2
   output [15:0] instruction;
   output wire inst_mem_err;
   output wire inst_mem_stall;
   output wire inst_mem_done;
   //output err; 
   
   // TODO: Your code here

   wire [15:0] pcNew;      //input of PC_reg
   wire [15:0] pcCurrent;  //output of PC_reg,
                           //intermediate value before adding 2

   //wire inst_mem_err;     //phase 2.1 align memory, if instruction memory has an error, disable the PC from incrementing
   //wire inst_mem_stall;   //phase 2.2 stall memory

   //Decision Order: stall > Halt > Halt
   //In my previous implementation, I use PCSrc as a second priority in pcNew MUX, 
   //which makes the stall generated by branch/jump_taken signal to be considered after the "Halt_fetch | normal stall"
   //Even though pcNew MUX has passed all the demo2 testing programs, this order may need to be reconsidered in the future demos
   //P.S. NOT SURE THE EXACT FUNCTION OF "Jump_IDEX" here...Need to reconsider in the future tests
   
   /*
   wire [15:0] branch_jump_pc_temp;
   reg16 branch_jump_flush_reg (.clk(clk), .rst(rst), .write(~inst_mem_stall), .wdata(branch_jump_pc), .rdata(branch_jump_pc_temp));
   
   assign pcNew = PCSrc                                                                   ?     branch_jump_pc_temp  : //branch_jump_pc_temp 
                  ~(Jump_IDEX) & (Halt_fetch | stall | inst_mem_err | inst_mem_stall)     ?     pcCurrent        : 
                                                                                                pcAdd2;
   */
   assign pcNew = PCSrc                                                   ?      branch_jump_pc  : //branch_jump_pc_temp 
                  ~(Jump_IDEX) & (Halt_fetch | stall | inst_mem_err )     ?      pcCurrent       : 
                                                                                 pcAdd2;

   
   //If Halt is after a jump, and Halt is decoded in Decode stage,
   //Meanwhile Jump is in Execute stage, need to prevent Halt_fetch stopping
   //PC from being updated, to succeed in jumping the PC

   wire [15:0] PC_addr_adder1_input_b;
   assign PC_addr_adder1_input_b = rst ? 16'h0000 : 16'h0002;
   cla_16b PC_addr_adder1(.sum(pcAdd2), .c_out(), .a(pcCurrent), .b(/*16'h0002*/PC_addr_adder1_input_b), .c_in(1'b0));        
   //c_out is overflow port, 
   //when there is an overflow error, an error will be output                               
   //err used to be output from c_out, but we no longer need err in demo2 testings


   reg16 PC_reg (.clk(clk), .rst(rst), .write(1'b1/*~rst*/), .wdata(pcNew/* & ~rst*/), .rdata(pcCurrent));

   /*
   memory2c Instruction_Memory(.data_out(instruction), .data_in(16'h0000), .addr(pcCurrent), 
   .enable(1'b1), .wr(1'b0), .createdump(1'b0), .clk(clk), .rst(rst)); //enable port is read enable
   */

   
   memory2c_align Instruction_Memory(
      .data_out(instruction), 
      .data_in(16'h0000), 
      .addr(pcCurrent), 
      .enable(~pcCurrent[0]),    //if ALU_out[0] is 1'b1, memory address is not aligned 
      .wr(1'b0), 
      .createdump(1'b0), 
      .clk(clk), 
      .rst(rst), 
      .err(inst_mem_err)
   );
   

   
   // stallmem Instruction_Memory(
   //    .DataOut(instruction), 
   //    .Done(inst_mem_done),                     //NOT SURE HOW TO CONNECT DONE SIGNAL
   //    .Stall(inst_mem_stall), 
   //    .CacheHit(), 
   //    .err(inst_mem_err), 
   //    .Addr(pcCurrent), 
   //    .DataIn(16'h0000), 
   //    .Rd(~pcCurrent[0]),     //enable port, if ALU_out[0] is 1'b1, memory address is not aligned
   //    .Wr(1'b0), 
   //    .createdump(1'b0), 
   //    .clk(clk), 
   //    .rst(rst)
   //    );

   
   
endmodule
