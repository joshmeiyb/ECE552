/*
   CS/ECE 552 Spring '20
  
   Filename        : wb.v
   Description     : This is the module for the overall Write Back stage of the processor.
*/
module wb (/* TODO: Add appropriate inputs/outputs for your WB stage here*/);

   // TODO: Your code here
   
endmodule
