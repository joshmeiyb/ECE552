/*
   CS/ECE 552 Spring '20
  
   Filename        : fetch.v
   Description     : This is the module for the overall fetch stage of the processor.
*/
module fetch (/* TODO: Add appropriate inputs/outputs for your fetch stage here*/);

   // TODO: Your code here
   
endmodule
