/*
   CS/ECE 552 Spring '20
  
   Filename        : fetch.v
   Description     : This is the module for the overall fetch stage of the processor.
*/
module fetch (clk, rst, /*err,*/ stall, 
               branch_jump_pc, PCSrc, Jump_IDEX,
               Halt_fetch, pcAdd2, 
               instruction
               );
   /* TODO: Add appropriate inputs/outputs for your fetch stage here*/
   
   input clk,rst;
   input stall;
   input [15:0] branch_jump_pc;  //used to be next_pc2
   input PCSrc;                  //branch_jump_taken signal
   input Jump_IDEX;
   input Halt_fetch;
   output [15:0] pcAdd2; //PC+2
   output [15:0] instruction;
   //output err; 
   
   // TODO: Your code here

   wire [15:0] pcNew;      //input of PC_reg
   wire [15:0] pcCurrent;  //output of PC_reg,
                           //intermediate value before adding 2

   //Decision Order: stall > Halt > Halt
   //In my previous implementation, I use PCSrc as a second priority in pcNew MUX, 
   //which makes the stall generated by branch/jump_taken signal to be considered after the "Halt_fetch | normal stall"
   //Even though pcNew MUX has passed all the demo2 testing programs, this order may need to be reconsidered in the future demos
   //P.S. NOT SURE THE EXACT FUNCTION OF "Jump_IDEX" here...Need to reconsider in the future tests
   assign pcNew = PCSrc                                  ?  branch_jump_pc   : 
                  ~(Jump_IDEX) & (Halt_fetch | stall)    ?  pcCurrent        : 
                                                            pcAdd2;
   //If Halt is after a jump, and Halt is decoded in Decode stage,
   //Meanwhile Jump is in Execute stage, need to prevent Halt_fetch stopping
   //PC from being updated, to succeed in jumping the PC

   wire [15:0] PC_addr_adder1_input_b;
   assign PC_addr_adder1_input_b = rst ? 16'h0000 : 16'h0002;
   cla_16b PC_addr_adder1(.sum(pcAdd2), .c_out(), .a(pcCurrent), .b(/*16'h0002*/PC_addr_adder1_input_b), .c_in(1'b0));        
   //c_out is overflow port, 
   //when there is an overflow error, an error will be output                               
   //err used to be output from c_out, but we no longer need err in demo2 testings


   reg16 PC_reg (.clk(clk), .rst(rst), .write(1'b1/*~rst*/), .wdata(pcNew/* & ~rst*/), .rdata(pcCurrent));

   memory2c Instruction_Memory(.data_out(instruction), .data_in(16'h0000), .addr(pcCurrent), 
   .enable(1'b1), .wr(1'b0), .createdump(1'b0), .clk(clk), .rst(rst)); //enable port is read enable

   
   
endmodule
