/*
    CS/ECE 552 Spring '22
    Homework #1, Problem 1

    1 input NOT
*/
module not1 (out, in1);
    output out;
    input in1;
    assign out = ~in1;
endmodule
